`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:32:44 11/08/2021 
// Design Name: 
// Module Name:    ScoreBoard 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ScoreBoard(
    input btn(3:0),
    input SW(7:0),
    input clk,
    output AN(3:0),
    output SEGMENT(7:0),
    output BTNX4
    );


endmodule
